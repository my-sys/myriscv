module riscv_soc(
	input	clock,
	input	reset,
);
  wire  core_clock; // @[riscv_soc.scala 42:20]
  wire  core_reset; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_aw_ready; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_aw_valid; // @[riscv_soc.scala 42:20]
  wire [63:0] core_io_axi_bus_aw_bits_awaddr; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_w_ready; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_w_valid; // @[riscv_soc.scala 42:20]
  wire [63:0] core_io_axi_bus_w_bits_wdata; // @[riscv_soc.scala 42:20]
  wire [7:0] core_io_axi_bus_w_bits_wstrb; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_w_bits_wlast; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_b_valid; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_ar_ready; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_ar_valid; // @[riscv_soc.scala 42:20]
  wire [63:0] core_io_axi_bus_ar_bits_araddr; // @[riscv_soc.scala 42:20]
  wire [7:0] core_io_axi_bus_ar_bits_arlen; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_r_valid; // @[riscv_soc.scala 42:20]
  wire [63:0] core_io_axi_bus_r_bits_rdata; // @[riscv_soc.scala 42:20]
  wire  core_io_axi_bus_r_bits_rlast; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram0_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram0_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram0_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram0_rdata; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram1_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram1_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram1_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram1_rdata; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram2_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram2_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram2_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram2_rdata; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram3_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram3_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram3_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram3_rdata; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram4_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram4_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram4_wmask; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram4_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram4_rdata; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram5_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram5_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram5_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram5_rdata; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram6_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram6_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram6_wmask; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram6_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram6_rdata; // @[riscv_soc.scala 42:20]
  wire [5:0] core_io_sram7_addr; // @[riscv_soc.scala 42:20]
  wire  core_io_sram7_wen; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram7_wdata; // @[riscv_soc.scala 42:20]
  wire [127:0] core_io_sram7_rdata; // @[riscv_soc.scala 42:20]
  wire  core_difftest_irq; // @[riscv_soc.scala 42:20]
  wire  core_difftest_peripheral; // @[riscv_soc.scala 42:20]
  wire  core_difftest_commit; // @[riscv_soc.scala 42:20]
  wire [63:0] core_difftest_pc; // @[riscv_soc.scala 42:20]
  wire [31:0] core_difftest_inst; // @[riscv_soc.scala 42:20]

  wire [63:0] core_inst_counter; // @[riscv_soc.scala 42:20]
  wire  axi_ram_clock; // @[riscv_soc.scala 43:23]
  wire  axi_ram_reset; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_aw_ready; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_aw_valid; // @[riscv_soc.scala 43:23]
  wire [63:0] axi_ram_io_ram_bus_aw_bits_awaddr; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_w_ready; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_w_valid; // @[riscv_soc.scala 43:23]
  wire [63:0] axi_ram_io_ram_bus_w_bits_wdata; // @[riscv_soc.scala 43:23]
  wire [7:0] axi_ram_io_ram_bus_w_bits_wstrb; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_w_bits_wlast; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_b_valid; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_ar_ready; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_ar_valid; // @[riscv_soc.scala 43:23]
  wire [63:0] axi_ram_io_ram_bus_ar_bits_araddr; // @[riscv_soc.scala 43:23]
  wire [7:0] axi_ram_io_ram_bus_ar_bits_arlen; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_r_valid; // @[riscv_soc.scala 43:23]
  wire [63:0] axi_ram_io_ram_bus_r_bits_rdata; // @[riscv_soc.scala 43:23]
  wire  axi_ram_io_ram_bus_r_bits_rlast; // @[riscv_soc.scala 43:23]
  wire  sram0_clock; // @[riscv_soc.scala 44:21]
  wire  sram0_reset; // @[riscv_soc.scala 44:21]
  wire [5:0] sram0_io_addr; // @[riscv_soc.scala 44:21]
  wire  sram0_io_wen; // @[riscv_soc.scala 44:21]
  wire [127:0] sram0_io_wmask; // @[riscv_soc.scala 44:21]
  wire [127:0] sram0_io_wdata; // @[riscv_soc.scala 44:21]
  wire [127:0] sram0_io_rdata; // @[riscv_soc.scala 44:21]
  wire  sram1_clock; // @[riscv_soc.scala 45:21]
  wire  sram1_reset; // @[riscv_soc.scala 45:21]
  wire [5:0] sram1_io_addr; // @[riscv_soc.scala 45:21]
  wire  sram1_io_wen; // @[riscv_soc.scala 45:21]
  wire [127:0] sram1_io_wmask; // @[riscv_soc.scala 45:21]
  wire [127:0] sram1_io_wdata; // @[riscv_soc.scala 45:21]
  wire [127:0] sram1_io_rdata; // @[riscv_soc.scala 45:21]
  wire  sram2_clock; // @[riscv_soc.scala 46:21]
  wire  sram2_reset; // @[riscv_soc.scala 46:21]
  wire [5:0] sram2_io_addr; // @[riscv_soc.scala 46:21]
  wire  sram2_io_wen; // @[riscv_soc.scala 46:21]
  wire [127:0] sram2_io_wmask; // @[riscv_soc.scala 46:21]
  wire [127:0] sram2_io_wdata; // @[riscv_soc.scala 46:21]
  wire [127:0] sram2_io_rdata; // @[riscv_soc.scala 46:21]
  wire  sram3_clock; // @[riscv_soc.scala 47:21]
  wire  sram3_reset; // @[riscv_soc.scala 47:21]
  wire [5:0] sram3_io_addr; // @[riscv_soc.scala 47:21]
  wire  sram3_io_wen; // @[riscv_soc.scala 47:21]
  wire [127:0] sram3_io_wmask; // @[riscv_soc.scala 47:21]
  wire [127:0] sram3_io_wdata; // @[riscv_soc.scala 47:21]
  wire [127:0] sram3_io_rdata; // @[riscv_soc.scala 47:21]
  wire  sram4_clock; // @[riscv_soc.scala 48:21]
  wire  sram4_reset; // @[riscv_soc.scala 48:21]
  wire [5:0] sram4_io_addr; // @[riscv_soc.scala 48:21]
  wire  sram4_io_wen; // @[riscv_soc.scala 48:21]
  wire [127:0] sram4_io_wmask; // @[riscv_soc.scala 48:21]
  wire [127:0] sram4_io_wdata; // @[riscv_soc.scala 48:21]
  wire [127:0] sram4_io_rdata; // @[riscv_soc.scala 48:21]
  wire  sram5_clock; // @[riscv_soc.scala 49:21]
  wire  sram5_reset; // @[riscv_soc.scala 49:21]
  wire [5:0] sram5_io_addr; // @[riscv_soc.scala 49:21]
  wire  sram5_io_wen; // @[riscv_soc.scala 49:21]
  wire [127:0] sram5_io_wmask; // @[riscv_soc.scala 49:21]
  wire [127:0] sram5_io_wdata; // @[riscv_soc.scala 49:21]
  wire [127:0] sram5_io_rdata; // @[riscv_soc.scala 49:21]
  wire  sram6_clock; // @[riscv_soc.scala 50:21]
  wire  sram6_reset; // @[riscv_soc.scala 50:21]
  wire [5:0] sram6_io_addr; // @[riscv_soc.scala 50:21]
  wire  sram6_io_wen; // @[riscv_soc.scala 50:21]
  wire [127:0] sram6_io_wmask; // @[riscv_soc.scala 50:21]
  wire [127:0] sram6_io_wdata; // @[riscv_soc.scala 50:21]
  wire [127:0] sram6_io_rdata; // @[riscv_soc.scala 50:21]
  wire  sram7_clock; // @[riscv_soc.scala 51:21]
  wire  sram7_reset; // @[riscv_soc.scala 51:21]
  wire [5:0] sram7_io_addr; // @[riscv_soc.scala 51:21]
  wire  sram7_io_wen; // @[riscv_soc.scala 51:21]
  wire [127:0] sram7_io_wmask; // @[riscv_soc.scala 51:21]
  wire [127:0] sram7_io_wdata; // @[riscv_soc.scala 51:21]
  wire [127:0] sram7_io_rdata; // @[riscv_soc.scala 51:21]
  wire [31:0] DIFFTEST_INST = core_difftest_inst;
  wire [63:0] difftest_inst = {{32'd0}, DIFFTEST_INST};
endmodule