module Decode(
  input         clock,
  input         reset,
  output        io_get_inst_ready,
  input         io_get_inst_valid,
  input  [31:0] io_get_inst_bits_inst,
  input  [63:0] io_get_inst_bits_pc,
  input         io_get_inst_bits_is_pre,
  output [4:0]  io_normal_rd_rs1_addr,
  input  [63:0] io_normal_rd_rs1_data,
  output [4:0]  io_normal_rd_rs2_addr,
  input  [63:0] io_normal_rd_rs2_data,
  output [11:0] io_csr_rd_csr_addr,
  input  [63:0] io_csr_rd_csr_data,
  input         io_op_datas_ready,
  output        io_op_datas_valid,
  output [2:0]  io_op_datas_bits_opType,
  output [6:0]  io_op_datas_bits_exuType,
  output [4:0]  io_op_datas_bits_rs1_addr,
  output [63:0] io_op_datas_bits_rs1_data,
  output [4:0]  io_op_datas_bits_rs2_addr,
  output [63:0] io_op_datas_bits_rs2_data,
  output [31:0] io_op_datas_bits_imm,
  output [63:0] io_op_datas_bits_pc,
  output [31:0] io_op_datas_bits_inst,
  output [4:0]  io_op_datas_bits_dest_addr,
  output        io_op_datas_bits_dest_is_reg,
  output        io_op_datas_bits_is_pre,
  output [11:0] io_op_datas_bits_csr_addr,
  output [63:0] io_op_datas_bits_csr_data,
  input         io_flush
);

  reg  reg_valid; // @[decode.scala 17:42]
  reg [2:0] reg_opType; // @[decode.scala 30:42]
  reg [6:0] reg_exuType; // @[decode.scala 31:42]
  reg [4:0] reg_rs1_addr; // @[decode.scala 32:42]
  reg [63:0] reg_rs1_data; // @[decode.scala 33:42]
  reg [4:0] reg_rs2_addr; // @[decode.scala 35:42]
  reg [63:0] reg_rs2_data; // @[decode.scala 36:42]
  reg [31:0] reg_imm; // @[decode.scala 37:42]
  reg [63:0] reg_pc; // @[decode.scala 38:50]
  reg [31:0] reg_inst; // @[decode.scala 40:42]
  reg [4:0] reg_dest_addr; // @[decode.scala 41:42]
  reg  reg_dest_is_reg; // @[decode.scala 42:38]
  reg [11:0] reg_csr_addr; // @[decode.scala 44:42]
  reg [63:0] reg_csr_data; // @[decode.scala 45:42]
  reg  reg_is_pre; // @[decode.scala 46:42]
  wire [4:0] rs2_addr = io_get_inst_bits_inst[24:20]; // @[decode.scala 54:35]
  wire [4:0] rs1_addr = io_get_inst_bits_inst[19:15]; // @[decode.scala 55:35]
  wire [11:0] csr_addr = io_get_inst_bits_inst[31:20]; // @[decode.scala 56:35]
  wire [4:0] dest_addr = io_get_inst_bits_inst[11:7]; // @[decode.scala 57:39]
  wire [2:0] fun = io_get_inst_bits_inst[14:12]; // @[decode.scala 59:23]
  wire [4:0] fun_exuType = {fun,io_get_inst_bits_inst[5],io_get_inst_bits_inst[3]}; // @[Cat.scala 33:92]
  wire [2:0] fun_op = {io_get_inst_bits_inst[6],io_get_inst_bits_inst[4],io_get_inst_bits_inst[2]}; // @[Cat.scala 33:92]
  wire  temp_system_is_pri = fun == 3'h0; // @[decode.scala 64:39]
  wire  temp_system_is_imm = io_get_inst_bits_inst[14]; // @[decode.scala 65:38]
  wire  temp_system_rs1 = temp_system_is_imm ? 1'h0 : 1'h1; // @[decode.scala 66:34]
  wire [6:0] _temp_system_T_1 = {io_get_inst_bits_inst[21:20],fun,io_get_inst_bits_inst[5],io_get_inst_bits_inst[3]}; // @[Cat.scala 33:92]
  wire [6:0] temp_system_1 = temp_system_is_pri ? _temp_system_T_1 : {{2'd0}, fun_exuType}; // @[decode.scala 70:53]
  wire [2:0] temp_system_2 = temp_system_is_pri ? 3'h0 : 3'h5; // @[decode.scala 71:12]
  wire  temp_system_3 = temp_system_is_pri ? 1'h0 : 1'h1; // @[decode.scala 71:72]
  wire  temp_system_4 = temp_system_is_pri ? 1'h0 : temp_system_rs1; // @[decode.scala 72:12]
  wire [3:0] temp_mem_itype = io_get_inst_bits_inst[5] ? 4'h3 : 4'hc; // @[decode.scala 73:33]
  wire  temp_mem_dest = io_get_inst_bits_inst[5] ? 1'h0 : 1'h1; // @[decode.scala 74:33]
  wire  temp_op_is_imm = ~io_get_inst_bits_inst[5]; // @[decode.scala 76:30]
  wire  is_sr = fun == 3'h5; // @[decode.scala 77:25]
  wire [5:0] temp_kk = {io_get_inst_bits_inst[30],fun,io_get_inst_bits_inst[5],io_get_inst_bits_inst[3]}; // @[Cat.scala 33:92]
  wire [5:0] _temp_op_exuType_T = is_sr ? temp_kk : {{1'd0}, fun_exuType}; // @[decode.scala 79:53]
  wire [5:0] temp_op_exuType = temp_op_is_imm ? _temp_op_exuType_T : temp_kk; // @[decode.scala 79:34]
  wire [3:0] _temp_op_itype_T_2 = fun == 3'h1 | is_sr ? 4'h4 : 4'hc; // @[decode.scala 80:51]
  wire [3:0] temp_op_itype = temp_op_is_imm ? _temp_op_itype_T_2 : 4'h6; // @[decode.scala 80:32]
  wire  temp_op_rs2 = temp_op_is_imm ? 1'h0 : 1'h1; // @[decode.scala 81:32]
  wire [2:0] _temp_op_T_1 = io_get_inst_bits_inst[25] ? 3'h5 : 3'h1; // @[decode.scala 82:60]
  wire [6:0] temp_jal_jalr_1 = io_get_inst_bits_inst[3] ? 7'h4e : 7'h4a; // @[decode.scala 86:12]
  wire [3:0] temp_jal_jalr_2 = io_get_inst_bits_inst[3] ? 4'h2 : 4'hc; // @[decode.scala 87:12]
  wire  temp_jal_jalr_4 = io_get_inst_bits_inst[3] ? 1'h0 : 1'h1; // @[decode.scala 88:12]
  wire [6:0] _T_1 = io_get_inst_bits_inst[5] ? 7'h0 : 7'h40; // @[decode.scala 91:59]
  wire [6:0] _T_2 = {2'h1,fun,io_get_inst_bits_inst[5],io_get_inst_bits_inst[3]}; // @[Cat.scala 33:92]
  wire [6:0] _T_3 = {2'h2,fun,io_get_inst_bits_inst[5],io_get_inst_bits_inst[3]}; // @[Cat.scala 33:92]
  wire  _T_5 = 3'h2 == fun_op; // @[Lookup.scala 31:38]
  wire  _T_7 = 3'h3 == fun_op; // @[Lookup.scala 31:38]
  wire  _T_9 = 3'h5 == fun_op; // @[Lookup.scala 31:38]
  wire  _T_11 = 3'h4 == fun_op; // @[Lookup.scala 31:38]
  wire  _T_13 = 3'h0 == fun_op; // @[Lookup.scala 31:38]
  wire  _T_15 = 3'h1 == fun_op; // @[Lookup.scala 31:38]
  wire  _T_17 = 3'h6 == fun_op; // @[Lookup.scala 31:38]
  wire [1:0] _T_18 = _T_17 ? 2'h3 : 2'h0; // @[Lookup.scala 34:39]
  wire [2:0] _T_19 = _T_15 ? 3'h4 : {{1'd0}, _T_18}; // @[Lookup.scala 34:39]
  wire [2:0] _T_20 = _T_13 ? 3'h0 : _T_19; // @[Lookup.scala 34:39]
  wire [2:0] _T_21 = _T_11 ? 3'h2 : _T_20; // @[Lookup.scala 34:39]
  wire [2:0] _T_22 = _T_9 ? 3'h2 : _T_21; // @[Lookup.scala 34:39]
  wire [6:0] _T_24 = _T_17 ? temp_system_1 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _T_25 = _T_15 ? _T_3 : _T_24; // @[Lookup.scala 34:39]
  wire [6:0] _T_26 = _T_13 ? {{2'd0}, fun_exuType} : _T_25; // @[Lookup.scala 34:39]
  wire [6:0] _T_27 = _T_11 ? _T_2 : _T_26; // @[Lookup.scala 34:39]
  wire [6:0] _T_28 = _T_9 ? temp_jal_jalr_1 : _T_27; // @[Lookup.scala 34:39]
  wire [2:0] _T_30 = _T_17 ? temp_system_2 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _T_31 = _T_15 ? 3'h0 : _T_30; // @[Lookup.scala 34:39]
  wire [3:0] _T_32 = _T_13 ? temp_mem_itype : {{1'd0}, _T_31}; // @[Lookup.scala 34:39]
  wire [3:0] _T_33 = _T_11 ? 4'h7 : _T_32; // @[Lookup.scala 34:39]
  wire [3:0] _T_34 = _T_9 ? temp_jal_jalr_2 : _T_33; // @[Lookup.scala 34:39]
  wire [3:0] _T_35 = _T_7 ? 4'h1 : _T_34; // @[Lookup.scala 34:39]
  wire [3:0] instType = _T_5 ? temp_op_itype : _T_35; // @[Lookup.scala 34:39]
  wire  _T_37 = _T_15 ? 1'h0 : _T_17 & temp_system_3; // @[Lookup.scala 34:39]
  wire  _T_38 = _T_13 ? temp_mem_dest : _T_37; // @[Lookup.scala 34:39]
  wire  _T_39 = _T_11 ? 1'h0 : _T_38; // @[Lookup.scala 34:39]
  wire  dest_is_reg = _T_5 | (_T_7 | (_T_9 | _T_39)); // @[Lookup.scala 34:39]
  wire  _T_43 = _T_15 ? 1'h0 : _T_17 & temp_system_4; // @[Lookup.scala 34:39]
  wire  _T_46 = _T_9 ? temp_jal_jalr_4 : _T_11 | (_T_13 | _T_43); // @[Lookup.scala 34:39]
  wire  _T_47 = _T_7 ? 1'h0 : _T_46; // @[Lookup.scala 34:39]
  wire  rs1_is_reg = _T_5 | _T_47; // @[Lookup.scala 34:39]
  wire  _T_52 = _T_9 ? 1'h0 : _T_11 | _T_13 & io_get_inst_bits_inst[5]; // @[Lookup.scala 34:39]
  wire  _T_53 = _T_7 ? 1'h0 : _T_52; // @[Lookup.scala 34:39]
  wire  rs2_is_reg = _T_5 ? temp_op_rs2 : _T_53; // @[Lookup.scala 34:39]
  wire [19:0] _imm_data_T_2 = io_get_inst_bits_inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _imm_data_T_4 = {_imm_data_T_2,csr_addr}; // @[Cat.scala 33:92]
  wire [31:0] _imm_data_T_6 = {io_get_inst_bits_inst[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [31:0] _imm_data_T_13 = {_imm_data_T_2,io_get_inst_bits_inst[31:25],dest_addr}; // @[Cat.scala 33:92]
  wire [11:0] _imm_data_T_16 = io_get_inst_bits_inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _imm_data_T_23 = {_imm_data_T_16,io_get_inst_bits_inst[19:12],io_get_inst_bits_inst[20],
    io_get_inst_bits_inst[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] _imm_data_T_33 = {_imm_data_T_2,io_get_inst_bits_inst[7],io_get_inst_bits_inst[30:25],
    io_get_inst_bits_inst[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] _imm_data_T_35 = {27'h0,rs1_addr}; // @[Cat.scala 33:92]
  wire [31:0] _imm_data_T_37 = {26'h0,io_get_inst_bits_inst[25:20]}; // @[Cat.scala 33:92]
  wire [31:0] _imm_data_T_39 = 4'hc == instType ? _imm_data_T_4 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _imm_data_T_41 = 4'h1 == instType ? _imm_data_T_6 : _imm_data_T_39; // @[Mux.scala 81:58]
  wire [31:0] _imm_data_T_43 = 4'h3 == instType ? _imm_data_T_13 : _imm_data_T_41; // @[Mux.scala 81:58]
  wire [31:0] _imm_data_T_45 = 4'h2 == instType ? _imm_data_T_23 : _imm_data_T_43; // @[Mux.scala 81:58]
  wire [31:0] _imm_data_T_47 = 4'h7 == instType ? _imm_data_T_33 : _imm_data_T_45; // @[Mux.scala 81:58]
  assign io_get_inst_ready = io_op_datas_ready; // @[decode.scala 21:31]
  assign io_normal_rd_rs1_addr = io_get_inst_bits_inst[19:15]; // @[decode.scala 55:35]
  assign io_normal_rd_rs2_addr = io_get_inst_bits_inst[24:20]; // @[decode.scala 54:35]
  assign io_csr_rd_csr_addr = io_get_inst_bits_inst[31:20]; // @[decode.scala 56:35]
  assign io_op_datas_valid = reg_valid; // @[decode.scala 161:57]
  assign io_op_datas_bits_opType = reg_opType; // @[decode.scala 146:49]
  assign io_op_datas_bits_exuType = reg_exuType; // @[decode.scala 147:49]
  assign io_op_datas_bits_rs1_addr = reg_rs1_addr; // @[decode.scala 148:49]
  assign io_op_datas_bits_rs1_data = reg_rs1_data; // @[decode.scala 149:49]
  assign io_op_datas_bits_rs2_addr = reg_rs2_addr; // @[decode.scala 150:49]
  assign io_op_datas_bits_rs2_data = reg_rs2_data; // @[decode.scala 151:49]
  assign io_op_datas_bits_imm = reg_imm; // @[decode.scala 152:49]
  assign io_op_datas_bits_pc = reg_pc; // @[decode.scala 153:57]
  assign io_op_datas_bits_inst = reg_inst; // @[decode.scala 154:49]
  assign io_op_datas_bits_dest_addr = reg_dest_addr; // @[decode.scala 155:49]
  assign io_op_datas_bits_dest_is_reg = reg_dest_is_reg; // @[decode.scala 156:41]
  assign io_op_datas_bits_is_pre = reg_is_pre; // @[decode.scala 160:49]
  assign io_op_datas_bits_csr_addr = reg_csr_addr; // @[decode.scala 158:49]
  assign io_op_datas_bits_csr_data = reg_csr_data; // @[decode.scala 159:49]
  always @(posedge clock) begin
    if (reset) begin // @[decode.scala 17:42]
      reg_valid <= 1'h0; // @[decode.scala 17:42]
    end else if (io_flush) begin // @[decode.scala 22:20]
      reg_valid <= 1'h0; // @[decode.scala 23:27]
    end else if (io_op_datas_ready) begin // @[decode.scala 25:28]
      reg_valid <= io_get_inst_valid; // @[decode.scala 26:41]
    end
    if (reset) begin // @[decode.scala 30:42]
      reg_opType <= 3'h0; // @[decode.scala 30:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      if (_T_5) begin // @[Lookup.scala 34:39]
        if (temp_op_is_imm) begin // @[decode.scala 82:26]
          reg_opType <= 3'h1;
        end else begin
          reg_opType <= _temp_op_T_1;
        end
      end else if (_T_7) begin // @[Lookup.scala 34:39]
        reg_opType <= 3'h1;
      end else begin
        reg_opType <= _T_22;
      end
    end
    if (reset) begin // @[decode.scala 31:42]
      reg_exuType <= 7'h0; // @[decode.scala 31:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      if (_T_5) begin // @[Lookup.scala 34:39]
        reg_exuType <= {{1'd0}, temp_op_exuType};
      end else if (_T_7) begin // @[Lookup.scala 34:39]
        reg_exuType <= _T_1;
      end else begin
        reg_exuType <= _T_28;
      end
    end
    if (reset) begin // @[decode.scala 32:42]
      reg_rs1_addr <= 5'h0; // @[decode.scala 32:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      if (rs1_is_reg) begin // @[decode.scala 116:34]
        reg_rs1_addr <= rs1_addr;
      end else begin
        reg_rs1_addr <= 5'h0;
      end
    end
    if (reset) begin // @[decode.scala 33:42]
      reg_rs1_data <= 64'h0; // @[decode.scala 33:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      if (rs1_is_reg) begin // @[decode.scala 117:34]
        reg_rs1_data <= io_normal_rd_rs1_data;
      end else begin
        reg_rs1_data <= 64'h0;
      end
    end
    if (reset) begin // @[decode.scala 35:42]
      reg_rs2_addr <= 5'h0; // @[decode.scala 35:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      if (rs2_is_reg) begin // @[decode.scala 118:34]
        reg_rs2_addr <= rs2_addr;
      end else begin
        reg_rs2_addr <= 5'h0;
      end
    end
    if (reset) begin // @[decode.scala 36:42]
      reg_rs2_data <= 64'h0; // @[decode.scala 36:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      if (rs2_is_reg) begin // @[decode.scala 119:34]
        reg_rs2_data <= io_normal_rd_rs2_data;
      end else begin
        reg_rs2_data <= 64'h0;
      end
    end
    if (reset) begin // @[decode.scala 37:42]
      reg_imm <= 32'h0; // @[decode.scala 37:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      if (4'h4 == instType) begin // @[Mux.scala 81:58]
        reg_imm <= _imm_data_T_37;
      end else if (4'h5 == instType) begin // @[Mux.scala 81:58]
        reg_imm <= _imm_data_T_35;
      end else begin
        reg_imm <= _imm_data_T_47;
      end
    end
    if (reset) begin // @[decode.scala 38:50]
      reg_pc <= 64'h0; // @[decode.scala 38:50]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      reg_pc <= io_get_inst_bits_pc; // @[decode.scala 131:41]
    end
    if (reset) begin // @[decode.scala 40:42]
      reg_inst <= 32'h0; // @[decode.scala 40:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      reg_inst <= io_get_inst_bits_inst; // @[decode.scala 133:41]
    end
    if (reset) begin // @[decode.scala 41:42]
      reg_dest_addr <= 5'h0; // @[decode.scala 41:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      reg_dest_addr <= dest_addr; // @[decode.scala 134:33]
    end
    if (reset) begin // @[decode.scala 42:38]
      reg_dest_is_reg <= 1'h0; // @[decode.scala 42:38]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      reg_dest_is_reg <= dest_is_reg; // @[decode.scala 135:33]
    end
    if (reset) begin // @[decode.scala 44:42]
      reg_csr_addr <= 12'h0; // @[decode.scala 44:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      reg_csr_addr <= csr_addr; // @[decode.scala 137:33]
    end
    if (reset) begin // @[decode.scala 45:42]
      reg_csr_data <= 64'h0; // @[decode.scala 45:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      reg_csr_data <= io_csr_rd_csr_data; // @[decode.scala 138:33]
    end
    if (reset) begin // @[decode.scala 46:42]
      reg_is_pre <= 1'h0; // @[decode.scala 46:42]
    end else if (io_op_datas_ready) begin // @[decode.scala 120:20]
      reg_is_pre <= io_get_inst_bits_is_pre; // @[decode.scala 139:41]
    end
  end
//   reg  reg_valid; // @[decode.scala 17:42]
//   reg [2:0] reg_opType; // @[decode.scala 30:42]
//   reg [6:0] reg_exuType; // @[decode.scala 31:42]
//   reg [4:0] reg_rs1_addr; // @[decode.scala 32:42]
//   reg [63:0] reg_rs1_data; // @[decode.scala 33:42]
//   reg [4:0] reg_rs2_addr; // @[decode.scala 35:42]
//   reg [63:0] reg_rs2_data; // @[decode.scala 36:42]
//   reg [31:0] reg_imm; // @[decode.scala 37:42]
//   reg [63:0] reg_pc; // @[decode.scala 38:50]
//   reg [31:0] reg_inst; // @[decode.scala 40:42]
//   reg [4:0] reg_dest_addr; // @[decode.scala 41:42]
//   reg  reg_dest_is_reg; // @[decode.scala 42:38]
//   reg [11:0] reg_csr_addr; // @[decode.scala 44:42]
//   reg [63:0] reg_csr_data; // @[decode.scala 45:42]
//   reg  reg_is_pre; // @[decode.scala 46:42]
//   wire [4:0] rs2_addr = io_get_inst_bits_inst[24:20]; // @[decode.scala 54:35]
//   wire [4:0] rs1_addr = io_get_inst_bits_inst[19:15]; // @[decode.scala 55:35]
//   wire [11:0] csr_addr = io_get_inst_bits_inst[31:20]; // @[decode.scala 56:35]
//   wire [4:0] dest_addr = io_get_inst_bits_inst[11:7]; // @[decode.scala 57:39]
//   wire [31:0] _T = io_get_inst_bits_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
//   wire  _T_1 = 32'h33 == _T; // @[Lookup.scala 31:38]
//   wire [31:0] _T_2 = io_get_inst_bits_inst & 32'h707f; // @[Lookup.scala 31:38]
//   wire  _T_3 = 32'h13 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_5 = 32'h1b == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_7 = 32'h3b == _T; // @[Lookup.scala 31:38]
//   wire  _T_9 = 32'h7033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_11 = 32'h7013 == _T_2; // @[Lookup.scala 31:38]
//   wire [31:0] _T_12 = io_get_inst_bits_inst & 32'h7f; // @[Lookup.scala 31:38]
//   wire  _T_13 = 32'h17 == _T_12; // @[Lookup.scala 31:38]
//   wire  _T_15 = 32'h63 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_17 = 32'h5063 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_19 = 32'h7063 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_21 = 32'h4063 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_23 = 32'h6063 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_25 = 32'h1063 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_27 = 32'h3073 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_29 = 32'h7073 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_31 = 32'h2073 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_33 = 32'h6073 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_35 = 32'h1073 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_37 = 32'h5073 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_39 = 32'h3003 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_41 = 32'h3 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_43 = 32'h4003 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_45 = 32'h1003 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_47 = 32'h5003 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_49 = 32'h37 == _T_12; // @[Lookup.scala 31:38]
//   wire  _T_51 = 32'h2003 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_53 = 32'h6003 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_55 = 32'h3023 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_57 = 32'h23 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_59 = 32'h1023 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_61 = 32'h1033 == _T; // @[Lookup.scala 31:38]
//   wire [31:0] _T_62 = io_get_inst_bits_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
//   wire  _T_63 = 32'h1013 == _T_62; // @[Lookup.scala 31:38]
//   wire  _T_65 = 32'h101b == _T; // @[Lookup.scala 31:38]
//   wire  _T_67 = 32'h103b == _T; // @[Lookup.scala 31:38]
//   wire  _T_69 = 32'h2033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_71 = 32'h2013 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_73 = 32'h3013 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_75 = 32'h3033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_77 = 32'h40005033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_79 = 32'h40005013 == _T_62; // @[Lookup.scala 31:38]
//   wire  _T_81 = 32'h4000501b == _T; // @[Lookup.scala 31:38]
//   wire  _T_83 = 32'h4000503b == _T; // @[Lookup.scala 31:38]
//   wire  _T_85 = 32'h5033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_87 = 32'h5013 == _T_62; // @[Lookup.scala 31:38]
//   wire  _T_89 = 32'h501b == _T; // @[Lookup.scala 31:38]
//   wire  _T_91 = 32'h503b == _T; // @[Lookup.scala 31:38]
//   wire  _T_93 = 32'h40000033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_95 = 32'h4000003b == _T; // @[Lookup.scala 31:38]
//   wire  _T_97 = 32'h2023 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_99 = 32'h6033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_101 = 32'h6013 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_103 = 32'h4033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_105 = 32'h4013 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_107 = 32'h2004033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_109 = 32'h2005033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_111 = 32'h200503b == _T; // @[Lookup.scala 31:38]
//   wire  _T_113 = 32'h200403b == _T; // @[Lookup.scala 31:38]
//   wire  _T_115 = 32'h2000033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_117 = 32'h2001033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_119 = 32'h2002033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_121 = 32'h2003033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_123 = 32'h200003b == _T; // @[Lookup.scala 31:38]
//   wire  _T_125 = 32'h2006033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_127 = 32'h2007033 == _T; // @[Lookup.scala 31:38]
//   wire  _T_129 = 32'h200703b == _T; // @[Lookup.scala 31:38]
//   wire  _T_131 = 32'h200603b == _T; // @[Lookup.scala 31:38]
//   wire  _T_133 = 32'h6f == _T_12; // @[Lookup.scala 31:38]
//   wire  _T_135 = 32'h67 == _T_2; // @[Lookup.scala 31:38]
//   wire  _T_137 = 32'h100073 == io_get_inst_bits_inst; // @[Lookup.scala 31:38]
//   wire  _T_139 = 32'h30200073 == io_get_inst_bits_inst; // @[Lookup.scala 31:38]
//   wire  _T_141 = 32'h73 == io_get_inst_bits_inst; // @[Lookup.scala 31:38]
//   wire  _T_143 = 32'h10200073 == io_get_inst_bits_inst; // @[Lookup.scala 31:38]
//   wire [31:0] _T_144 = io_get_inst_bits_inst & 32'hf00fffff; // @[Lookup.scala 31:38]
//   wire  _T_145 = 32'hf == _T_144; // @[Lookup.scala 31:38]
//   wire  _T_147 = 32'h100f == io_get_inst_bits_inst; // @[Lookup.scala 31:38]
//   wire [31:0] _T_148 = io_get_inst_bits_inst & 32'hfe007fff; // @[Lookup.scala 31:38]
//   wire  _T_149 = 32'h12000073 == _T_148; // @[Lookup.scala 31:38]
//   wire [2:0] _T_150 = _T_149 ? 3'h6 : 3'h0; // @[Lookup.scala 34:39]
//   wire [2:0] _T_151 = _T_147 ? 3'h6 : _T_150; // @[Lookup.scala 34:39]
//   wire [2:0] _T_152 = _T_145 ? 3'h6 : _T_151; // @[Lookup.scala 34:39]
//   wire [2:0] _T_153 = _T_143 ? 3'h4 : _T_152; // @[Lookup.scala 34:39]
//   wire [2:0] _T_154 = _T_141 ? 3'h4 : _T_153; // @[Lookup.scala 34:39]
//   wire [2:0] _T_155 = _T_139 ? 3'h4 : _T_154; // @[Lookup.scala 34:39]
//   wire [2:0] _T_156 = _T_137 ? 3'h4 : _T_155; // @[Lookup.scala 34:39]
//   wire [2:0] _T_157 = _T_135 ? 3'h1 : _T_156; // @[Lookup.scala 34:39]
//   wire [2:0] _T_158 = _T_133 ? 3'h1 : _T_157; // @[Lookup.scala 34:39]
//   wire [2:0] _T_159 = _T_131 ? 3'h3 : _T_158; // @[Lookup.scala 34:39]
//   wire [2:0] _T_160 = _T_129 ? 3'h3 : _T_159; // @[Lookup.scala 34:39]
//   wire [2:0] _T_161 = _T_127 ? 3'h3 : _T_160; // @[Lookup.scala 34:39]
//   wire [2:0] _T_162 = _T_125 ? 3'h3 : _T_161; // @[Lookup.scala 34:39]
//   wire [2:0] _T_163 = _T_123 ? 3'h3 : _T_162; // @[Lookup.scala 34:39]
//   wire [2:0] _T_164 = _T_121 ? 3'h3 : _T_163; // @[Lookup.scala 34:39]
//   wire [2:0] _T_165 = _T_119 ? 3'h3 : _T_164; // @[Lookup.scala 34:39]
//   wire [2:0] _T_166 = _T_117 ? 3'h3 : _T_165; // @[Lookup.scala 34:39]
//   wire [2:0] _T_167 = _T_115 ? 3'h3 : _T_166; // @[Lookup.scala 34:39]
//   wire [2:0] _T_168 = _T_113 ? 3'h3 : _T_167; // @[Lookup.scala 34:39]
//   wire [2:0] _T_169 = _T_111 ? 3'h3 : _T_168; // @[Lookup.scala 34:39]
//   wire [2:0] _T_170 = _T_109 ? 3'h3 : _T_169; // @[Lookup.scala 34:39]
//   wire [2:0] _T_171 = _T_107 ? 3'h3 : _T_170; // @[Lookup.scala 34:39]
//   wire [2:0] _T_172 = _T_105 ? 3'h2 : _T_171; // @[Lookup.scala 34:39]
//   wire [2:0] _T_173 = _T_103 ? 3'h2 : _T_172; // @[Lookup.scala 34:39]
//   wire [2:0] _T_174 = _T_101 ? 3'h2 : _T_173; // @[Lookup.scala 34:39]
//   wire [2:0] _T_175 = _T_99 ? 3'h2 : _T_174; // @[Lookup.scala 34:39]
//   wire [2:0] _T_176 = _T_97 ? 3'h5 : _T_175; // @[Lookup.scala 34:39]
//   wire [2:0] _T_177 = _T_95 ? 3'h2 : _T_176; // @[Lookup.scala 34:39]
//   wire [2:0] _T_178 = _T_93 ? 3'h2 : _T_177; // @[Lookup.scala 34:39]
//   wire [2:0] _T_179 = _T_91 ? 3'h2 : _T_178; // @[Lookup.scala 34:39]
//   wire [2:0] _T_180 = _T_89 ? 3'h2 : _T_179; // @[Lookup.scala 34:39]
//   wire [2:0] _T_181 = _T_87 ? 3'h2 : _T_180; // @[Lookup.scala 34:39]
//   wire [2:0] _T_182 = _T_85 ? 3'h2 : _T_181; // @[Lookup.scala 34:39]
//   wire [2:0] _T_183 = _T_83 ? 3'h2 : _T_182; // @[Lookup.scala 34:39]
//   wire [2:0] _T_184 = _T_81 ? 3'h2 : _T_183; // @[Lookup.scala 34:39]
//   wire [2:0] _T_185 = _T_79 ? 3'h2 : _T_184; // @[Lookup.scala 34:39]
//   wire [2:0] _T_186 = _T_77 ? 3'h2 : _T_185; // @[Lookup.scala 34:39]
//   wire [2:0] _T_187 = _T_75 ? 3'h2 : _T_186; // @[Lookup.scala 34:39]
//   wire [2:0] _T_188 = _T_73 ? 3'h2 : _T_187; // @[Lookup.scala 34:39]
//   wire [2:0] _T_189 = _T_71 ? 3'h2 : _T_188; // @[Lookup.scala 34:39]
//   wire [2:0] _T_190 = _T_69 ? 3'h2 : _T_189; // @[Lookup.scala 34:39]
//   wire [2:0] _T_191 = _T_67 ? 3'h2 : _T_190; // @[Lookup.scala 34:39]
//   wire [2:0] _T_192 = _T_65 ? 3'h2 : _T_191; // @[Lookup.scala 34:39]
//   wire [2:0] _T_193 = _T_63 ? 3'h2 : _T_192; // @[Lookup.scala 34:39]
//   wire [2:0] _T_194 = _T_61 ? 3'h2 : _T_193; // @[Lookup.scala 34:39]
//   wire [2:0] _T_195 = _T_59 ? 3'h5 : _T_194; // @[Lookup.scala 34:39]
//   wire [2:0] _T_196 = _T_57 ? 3'h5 : _T_195; // @[Lookup.scala 34:39]
//   wire [2:0] _T_197 = _T_55 ? 3'h5 : _T_196; // @[Lookup.scala 34:39]
//   wire [2:0] _T_198 = _T_53 ? 3'h5 : _T_197; // @[Lookup.scala 34:39]
//   wire [2:0] _T_199 = _T_51 ? 3'h5 : _T_198; // @[Lookup.scala 34:39]
//   wire [2:0] _T_200 = _T_49 ? 3'h2 : _T_199; // @[Lookup.scala 34:39]
//   wire [2:0] _T_201 = _T_47 ? 3'h5 : _T_200; // @[Lookup.scala 34:39]
//   wire [2:0] _T_202 = _T_45 ? 3'h5 : _T_201; // @[Lookup.scala 34:39]
//   wire [2:0] _T_203 = _T_43 ? 3'h5 : _T_202; // @[Lookup.scala 34:39]
//   wire [2:0] _T_204 = _T_41 ? 3'h5 : _T_203; // @[Lookup.scala 34:39]
//   wire [2:0] _T_205 = _T_39 ? 3'h5 : _T_204; // @[Lookup.scala 34:39]
//   wire [2:0] _T_206 = _T_37 ? 3'h4 : _T_205; // @[Lookup.scala 34:39]
//   wire [2:0] _T_207 = _T_35 ? 3'h4 : _T_206; // @[Lookup.scala 34:39]
//   wire [2:0] _T_208 = _T_33 ? 3'h4 : _T_207; // @[Lookup.scala 34:39]
//   wire [2:0] _T_209 = _T_31 ? 3'h4 : _T_208; // @[Lookup.scala 34:39]
//   wire [2:0] _T_210 = _T_29 ? 3'h4 : _T_209; // @[Lookup.scala 34:39]
//   wire [2:0] _T_211 = _T_27 ? 3'h4 : _T_210; // @[Lookup.scala 34:39]
//   wire [2:0] _T_212 = _T_25 ? 3'h1 : _T_211; // @[Lookup.scala 34:39]
//   wire [2:0] _T_213 = _T_23 ? 3'h1 : _T_212; // @[Lookup.scala 34:39]
//   wire [2:0] _T_214 = _T_21 ? 3'h1 : _T_213; // @[Lookup.scala 34:39]
//   wire [2:0] _T_215 = _T_19 ? 3'h1 : _T_214; // @[Lookup.scala 34:39]
//   wire [2:0] _T_216 = _T_17 ? 3'h1 : _T_215; // @[Lookup.scala 34:39]
//   wire [2:0] _T_217 = _T_15 ? 3'h1 : _T_216; // @[Lookup.scala 34:39]
//   wire [2:0] _T_218 = _T_13 ? 3'h2 : _T_217; // @[Lookup.scala 34:39]
//   wire [2:0] _T_219 = _T_11 ? 3'h2 : _T_218; // @[Lookup.scala 34:39]
//   wire [2:0] _T_220 = _T_9 ? 3'h2 : _T_219; // @[Lookup.scala 34:39]
//   wire [2:0] _T_221 = _T_7 ? 3'h2 : _T_220; // @[Lookup.scala 34:39]
//   wire [2:0] _T_222 = _T_5 ? 3'h2 : _T_221; // @[Lookup.scala 34:39]
//   wire [1:0] _T_224 = _T_149 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
//   wire [2:0] _T_225 = _T_147 ? 3'h5 : {{1'd0}, _T_224}; // @[Lookup.scala 34:39]
//   wire [2:0] _T_226 = _T_145 ? 3'h1 : _T_225; // @[Lookup.scala 34:39]
//   wire [6:0] _T_227 = _T_143 ? 7'h62 : {{4'd0}, _T_226}; // @[Lookup.scala 34:39]
//   wire [6:0] _T_228 = _T_141 ? 7'h2 : _T_227; // @[Lookup.scala 34:39]
//   wire [6:0] _T_229 = _T_139 ? 7'h42 : _T_228; // @[Lookup.scala 34:39]
//   wire [6:0] _T_230 = _T_137 ? 7'h22 : _T_229; // @[Lookup.scala 34:39]
//   wire [6:0] _T_231 = _T_135 ? 7'ha : _T_230; // @[Lookup.scala 34:39]
//   wire [6:0] _T_232 = _T_133 ? 7'he : _T_231; // @[Lookup.scala 34:39]
//   wire [6:0] _T_233 = _T_131 ? 7'h1b : _T_232; // @[Lookup.scala 34:39]
//   wire [6:0] _T_234 = _T_129 ? 7'h1f : _T_233; // @[Lookup.scala 34:39]
//   wire [6:0] _T_235 = _T_127 ? 7'h1e : _T_234; // @[Lookup.scala 34:39]
//   wire [6:0] _T_236 = _T_125 ? 7'h1a : _T_235; // @[Lookup.scala 34:39]
//   wire [6:0] _T_237 = _T_123 ? 7'h3 : _T_236; // @[Lookup.scala 34:39]
//   wire [6:0] _T_238 = _T_121 ? 7'he : _T_237; // @[Lookup.scala 34:39]
//   wire [6:0] _T_239 = _T_119 ? 7'ha : _T_238; // @[Lookup.scala 34:39]
//   wire [6:0] _T_240 = _T_117 ? 7'h6 : _T_239; // @[Lookup.scala 34:39]
//   wire [6:0] _T_241 = _T_115 ? 7'h2 : _T_240; // @[Lookup.scala 34:39]
//   wire [6:0] _T_242 = _T_113 ? 7'h13 : _T_241; // @[Lookup.scala 34:39]
//   wire [6:0] _T_243 = _T_111 ? 7'h17 : _T_242; // @[Lookup.scala 34:39]
//   wire [6:0] _T_244 = _T_109 ? 7'h16 : _T_243; // @[Lookup.scala 34:39]
//   wire [6:0] _T_245 = _T_107 ? 7'h12 : _T_244; // @[Lookup.scala 34:39]
//   wire [6:0] _T_246 = _T_105 ? 7'h10 : _T_245; // @[Lookup.scala 34:39]
//   wire [6:0] _T_247 = _T_103 ? 7'h12 : _T_246; // @[Lookup.scala 34:39]
//   wire [6:0] _T_248 = _T_101 ? 7'h18 : _T_247; // @[Lookup.scala 34:39]
//   wire [6:0] _T_249 = _T_99 ? 7'h1a : _T_248; // @[Lookup.scala 34:39]
//   wire [6:0] _T_250 = _T_97 ? 7'ha : _T_249; // @[Lookup.scala 34:39]
//   wire [6:0] _T_251 = _T_95 ? 7'h23 : _T_250; // @[Lookup.scala 34:39]
//   wire [6:0] _T_252 = _T_93 ? 7'h22 : _T_251; // @[Lookup.scala 34:39]
//   wire [6:0] _T_253 = _T_91 ? 7'h17 : _T_252; // @[Lookup.scala 34:39]
//   wire [6:0] _T_254 = _T_89 ? 7'h15 : _T_253; // @[Lookup.scala 34:39]
//   wire [6:0] _T_255 = _T_87 ? 7'h14 : _T_254; // @[Lookup.scala 34:39]
//   wire [6:0] _T_256 = _T_85 ? 7'h16 : _T_255; // @[Lookup.scala 34:39]
//   wire [6:0] _T_257 = _T_83 ? 7'h37 : _T_256; // @[Lookup.scala 34:39]
//   wire [6:0] _T_258 = _T_81 ? 7'h35 : _T_257; // @[Lookup.scala 34:39]
//   wire [6:0] _T_259 = _T_79 ? 7'h34 : _T_258; // @[Lookup.scala 34:39]
//   wire [6:0] _T_260 = _T_77 ? 7'h36 : _T_259; // @[Lookup.scala 34:39]
//   wire [6:0] _T_261 = _T_75 ? 7'h2e : _T_260; // @[Lookup.scala 34:39]
//   wire [6:0] _T_262 = _T_73 ? 7'h2c : _T_261; // @[Lookup.scala 34:39]
//   wire [6:0] _T_263 = _T_71 ? 7'h28 : _T_262; // @[Lookup.scala 34:39]
//   wire [6:0] _T_264 = _T_69 ? 7'h2a : _T_263; // @[Lookup.scala 34:39]
//   wire [6:0] _T_265 = _T_67 ? 7'h7 : _T_264; // @[Lookup.scala 34:39]
//   wire [6:0] _T_266 = _T_65 ? 7'h5 : _T_265; // @[Lookup.scala 34:39]
//   wire [6:0] _T_267 = _T_63 ? 7'h4 : _T_266; // @[Lookup.scala 34:39]
//   wire [6:0] _T_268 = _T_61 ? 7'h6 : _T_267; // @[Lookup.scala 34:39]
//   wire [6:0] _T_269 = _T_59 ? 7'h6 : _T_268; // @[Lookup.scala 34:39]
//   wire [6:0] _T_270 = _T_57 ? 7'h2 : _T_269; // @[Lookup.scala 34:39]
//   wire [6:0] _T_271 = _T_55 ? 7'he : _T_270; // @[Lookup.scala 34:39]
//   wire [6:0] _T_272 = _T_53 ? 7'h18 : _T_271; // @[Lookup.scala 34:39]
//   wire [6:0] _T_273 = _T_51 ? 7'h8 : _T_272; // @[Lookup.scala 34:39]
//   wire [6:0] _T_274 = _T_49 ? 7'h40 : _T_273; // @[Lookup.scala 34:39]
//   wire [6:0] _T_275 = _T_47 ? 7'h14 : _T_274; // @[Lookup.scala 34:39]
//   wire [6:0] _T_276 = _T_45 ? 7'h4 : _T_275; // @[Lookup.scala 34:39]
//   wire [6:0] _T_277 = _T_43 ? 7'h10 : _T_276; // @[Lookup.scala 34:39]
//   wire [6:0] _T_278 = _T_41 ? 7'h0 : _T_277; // @[Lookup.scala 34:39]
//   wire [6:0] _T_279 = _T_39 ? 7'hc : _T_278; // @[Lookup.scala 34:39]
//   wire [6:0] _T_280 = _T_37 ? 7'h16 : _T_279; // @[Lookup.scala 34:39]
//   wire [6:0] _T_281 = _T_35 ? 7'h6 : _T_280; // @[Lookup.scala 34:39]
//   wire [6:0] _T_282 = _T_33 ? 7'h1a : _T_281; // @[Lookup.scala 34:39]
//   wire [6:0] _T_283 = _T_31 ? 7'ha : _T_282; // @[Lookup.scala 34:39]
//   wire [6:0] _T_284 = _T_29 ? 7'h1e : _T_283; // @[Lookup.scala 34:39]
//   wire [6:0] _T_285 = _T_27 ? 7'he : _T_284; // @[Lookup.scala 34:39]
//   wire [6:0] _T_286 = _T_25 ? 7'h26 : _T_285; // @[Lookup.scala 34:39]
//   wire [6:0] _T_287 = _T_23 ? 7'h3a : _T_286; // @[Lookup.scala 34:39]
//   wire [6:0] _T_288 = _T_21 ? 7'h32 : _T_287; // @[Lookup.scala 34:39]
//   wire [6:0] _T_289 = _T_19 ? 7'h3e : _T_288; // @[Lookup.scala 34:39]
//   wire [6:0] _T_290 = _T_17 ? 7'h36 : _T_289; // @[Lookup.scala 34:39]
//   wire [6:0] _T_291 = _T_15 ? 7'h22 : _T_290; // @[Lookup.scala 34:39]
//   wire [6:0] _T_292 = _T_13 ? 7'h60 : _T_291; // @[Lookup.scala 34:39]
//   wire [6:0] _T_293 = _T_11 ? 7'h1c : _T_292; // @[Lookup.scala 34:39]
//   wire [6:0] _T_294 = _T_9 ? 7'h1e : _T_293; // @[Lookup.scala 34:39]
//   wire [6:0] _T_295 = _T_7 ? 7'h3 : _T_294; // @[Lookup.scala 34:39]
//   wire [6:0] _T_296 = _T_5 ? 7'h1 : _T_295; // @[Lookup.scala 34:39]
//   wire [3:0] _T_305 = _T_135 ? 4'hc : 4'h0; // @[Lookup.scala 34:39]
//   wire [3:0] _T_306 = _T_133 ? 4'h2 : _T_305; // @[Lookup.scala 34:39]
//   wire [3:0] _T_307 = _T_131 ? 4'h6 : _T_306; // @[Lookup.scala 34:39]
//   wire [3:0] _T_308 = _T_129 ? 4'h6 : _T_307; // @[Lookup.scala 34:39]
//   wire [3:0] _T_309 = _T_127 ? 4'h6 : _T_308; // @[Lookup.scala 34:39]
//   wire [3:0] _T_310 = _T_125 ? 4'h6 : _T_309; // @[Lookup.scala 34:39]
//   wire [3:0] _T_311 = _T_123 ? 4'h6 : _T_310; // @[Lookup.scala 34:39]
//   wire [3:0] _T_312 = _T_121 ? 4'h6 : _T_311; // @[Lookup.scala 34:39]
//   wire [3:0] _T_313 = _T_119 ? 4'h6 : _T_312; // @[Lookup.scala 34:39]
//   wire [3:0] _T_314 = _T_117 ? 4'h6 : _T_313; // @[Lookup.scala 34:39]
//   wire [3:0] _T_315 = _T_115 ? 4'h6 : _T_314; // @[Lookup.scala 34:39]
//   wire [3:0] _T_316 = _T_113 ? 4'h6 : _T_315; // @[Lookup.scala 34:39]
//   wire [3:0] _T_317 = _T_111 ? 4'h6 : _T_316; // @[Lookup.scala 34:39]
//   wire [3:0] _T_318 = _T_109 ? 4'h6 : _T_317; // @[Lookup.scala 34:39]
//   wire [3:0] _T_319 = _T_107 ? 4'h6 : _T_318; // @[Lookup.scala 34:39]
//   wire [3:0] _T_320 = _T_105 ? 4'hc : _T_319; // @[Lookup.scala 34:39]
//   wire [3:0] _T_321 = _T_103 ? 4'h6 : _T_320; // @[Lookup.scala 34:39]
//   wire [3:0] _T_322 = _T_101 ? 4'hc : _T_321; // @[Lookup.scala 34:39]
//   wire [3:0] _T_323 = _T_99 ? 4'h6 : _T_322; // @[Lookup.scala 34:39]
//   wire [3:0] _T_324 = _T_97 ? 4'h3 : _T_323; // @[Lookup.scala 34:39]
//   wire [3:0] _T_325 = _T_95 ? 4'h6 : _T_324; // @[Lookup.scala 34:39]
//   wire [3:0] _T_326 = _T_93 ? 4'h6 : _T_325; // @[Lookup.scala 34:39]
//   wire [3:0] _T_327 = _T_91 ? 4'h6 : _T_326; // @[Lookup.scala 34:39]
//   wire [3:0] _T_328 = _T_89 ? 4'h4 : _T_327; // @[Lookup.scala 34:39]
//   wire [3:0] _T_329 = _T_87 ? 4'h4 : _T_328; // @[Lookup.scala 34:39]
//   wire [3:0] _T_330 = _T_85 ? 4'h6 : _T_329; // @[Lookup.scala 34:39]
//   wire [3:0] _T_331 = _T_83 ? 4'h6 : _T_330; // @[Lookup.scala 34:39]
//   wire [3:0] _T_332 = _T_81 ? 4'h4 : _T_331; // @[Lookup.scala 34:39]
//   wire [3:0] _T_333 = _T_79 ? 4'h4 : _T_332; // @[Lookup.scala 34:39]
//   wire [3:0] _T_334 = _T_77 ? 4'h6 : _T_333; // @[Lookup.scala 34:39]
//   wire [3:0] _T_335 = _T_75 ? 4'h6 : _T_334; // @[Lookup.scala 34:39]
//   wire [3:0] _T_336 = _T_73 ? 4'hc : _T_335; // @[Lookup.scala 34:39]
//   wire [3:0] _T_337 = _T_71 ? 4'hc : _T_336; // @[Lookup.scala 34:39]
//   wire [3:0] _T_338 = _T_69 ? 4'h6 : _T_337; // @[Lookup.scala 34:39]
//   wire [3:0] _T_339 = _T_67 ? 4'h6 : _T_338; // @[Lookup.scala 34:39]
//   wire [3:0] _T_340 = _T_65 ? 4'h4 : _T_339; // @[Lookup.scala 34:39]
//   wire [3:0] _T_341 = _T_63 ? 4'h4 : _T_340; // @[Lookup.scala 34:39]
//   wire [3:0] _T_342 = _T_61 ? 4'h6 : _T_341; // @[Lookup.scala 34:39]
//   wire [3:0] _T_343 = _T_59 ? 4'h3 : _T_342; // @[Lookup.scala 34:39]
//   wire [3:0] _T_344 = _T_57 ? 4'h3 : _T_343; // @[Lookup.scala 34:39]
//   wire [3:0] _T_345 = _T_55 ? 4'h3 : _T_344; // @[Lookup.scala 34:39]
//   wire [3:0] _T_346 = _T_53 ? 4'hc : _T_345; // @[Lookup.scala 34:39]
//   wire [3:0] _T_347 = _T_51 ? 4'hc : _T_346; // @[Lookup.scala 34:39]
//   wire [3:0] _T_348 = _T_49 ? 4'h1 : _T_347; // @[Lookup.scala 34:39]
//   wire [3:0] _T_349 = _T_47 ? 4'hc : _T_348; // @[Lookup.scala 34:39]
//   wire [3:0] _T_350 = _T_45 ? 4'hc : _T_349; // @[Lookup.scala 34:39]
//   wire [3:0] _T_351 = _T_43 ? 4'hc : _T_350; // @[Lookup.scala 34:39]
//   wire [3:0] _T_352 = _T_41 ? 4'hc : _T_351; // @[Lookup.scala 34:39]
//   wire [3:0] _T_353 = _T_39 ? 4'hc : _T_352; // @[Lookup.scala 34:39]
//   wire [3:0] _T_354 = _T_37 ? 4'h5 : _T_353; // @[Lookup.scala 34:39]
//   wire [3:0] _T_355 = _T_35 ? 4'h5 : _T_354; // @[Lookup.scala 34:39]
//   wire [3:0] _T_356 = _T_33 ? 4'h5 : _T_355; // @[Lookup.scala 34:39]
//   wire [3:0] _T_357 = _T_31 ? 4'h5 : _T_356; // @[Lookup.scala 34:39]
//   wire [3:0] _T_358 = _T_29 ? 4'h5 : _T_357; // @[Lookup.scala 34:39]
//   wire [3:0] _T_359 = _T_27 ? 4'h5 : _T_358; // @[Lookup.scala 34:39]
//   wire [3:0] _T_360 = _T_25 ? 4'h7 : _T_359; // @[Lookup.scala 34:39]
//   wire [3:0] _T_361 = _T_23 ? 4'h7 : _T_360; // @[Lookup.scala 34:39]
//   wire [3:0] _T_362 = _T_21 ? 4'h7 : _T_361; // @[Lookup.scala 34:39]
//   wire [3:0] _T_363 = _T_19 ? 4'h7 : _T_362; // @[Lookup.scala 34:39]
//   wire [3:0] _T_364 = _T_17 ? 4'h7 : _T_363; // @[Lookup.scala 34:39]
//   wire [3:0] _T_365 = _T_15 ? 4'h7 : _T_364; // @[Lookup.scala 34:39]
//   wire [3:0] _T_366 = _T_13 ? 4'h1 : _T_365; // @[Lookup.scala 34:39]
//   wire [3:0] _T_367 = _T_11 ? 4'hc : _T_366; // @[Lookup.scala 34:39]
//   wire [3:0] _T_368 = _T_9 ? 4'h6 : _T_367; // @[Lookup.scala 34:39]
//   wire [3:0] _T_369 = _T_7 ? 4'h6 : _T_368; // @[Lookup.scala 34:39]
//   wire [3:0] _T_370 = _T_5 ? 4'hc : _T_369; // @[Lookup.scala 34:39]
//   wire [3:0] _T_371 = _T_3 ? 4'hc : _T_370; // @[Lookup.scala 34:39]
//   wire [3:0] instType = _T_1 ? 4'h6 : _T_371; // @[Lookup.scala 34:39]
//   wire [1:0] _T_379 = _T_135 ? 2'h1 : 2'h0; // @[Lookup.scala 34:39]
//   wire [1:0] _T_380 = _T_133 ? 2'h1 : _T_379; // @[Lookup.scala 34:39]
//   wire [1:0] _T_381 = _T_131 ? 2'h1 : _T_380; // @[Lookup.scala 34:39]
//   wire [1:0] _T_382 = _T_129 ? 2'h1 : _T_381; // @[Lookup.scala 34:39]
//   wire [1:0] _T_383 = _T_127 ? 2'h1 : _T_382; // @[Lookup.scala 34:39]
//   wire [1:0] _T_384 = _T_125 ? 2'h1 : _T_383; // @[Lookup.scala 34:39]
//   wire [1:0] _T_385 = _T_123 ? 2'h1 : _T_384; // @[Lookup.scala 34:39]
//   wire [1:0] _T_386 = _T_121 ? 2'h1 : _T_385; // @[Lookup.scala 34:39]
//   wire [1:0] _T_387 = _T_119 ? 2'h1 : _T_386; // @[Lookup.scala 34:39]
//   wire [1:0] _T_388 = _T_117 ? 2'h1 : _T_387; // @[Lookup.scala 34:39]
//   wire [1:0] _T_389 = _T_115 ? 2'h1 : _T_388; // @[Lookup.scala 34:39]
//   wire [1:0] _T_390 = _T_113 ? 2'h1 : _T_389; // @[Lookup.scala 34:39]
//   wire [1:0] _T_391 = _T_111 ? 2'h1 : _T_390; // @[Lookup.scala 34:39]
//   wire [1:0] _T_392 = _T_109 ? 2'h1 : _T_391; // @[Lookup.scala 34:39]
//   wire [1:0] _T_393 = _T_107 ? 2'h1 : _T_392; // @[Lookup.scala 34:39]
//   wire [1:0] _T_394 = _T_105 ? 2'h1 : _T_393; // @[Lookup.scala 34:39]
//   wire [1:0] _T_395 = _T_103 ? 2'h1 : _T_394; // @[Lookup.scala 34:39]
//   wire [1:0] _T_396 = _T_101 ? 2'h1 : _T_395; // @[Lookup.scala 34:39]
//   wire [1:0] _T_397 = _T_99 ? 2'h1 : _T_396; // @[Lookup.scala 34:39]
//   wire [1:0] _T_398 = _T_97 ? 2'h0 : _T_397; // @[Lookup.scala 34:39]
//   wire [1:0] _T_399 = _T_95 ? 2'h1 : _T_398; // @[Lookup.scala 34:39]
//   wire [1:0] _T_400 = _T_93 ? 2'h1 : _T_399; // @[Lookup.scala 34:39]
//   wire [1:0] _T_401 = _T_91 ? 2'h1 : _T_400; // @[Lookup.scala 34:39]
//   wire [1:0] _T_402 = _T_89 ? 2'h1 : _T_401; // @[Lookup.scala 34:39]
//   wire [1:0] _T_403 = _T_87 ? 2'h1 : _T_402; // @[Lookup.scala 34:39]
//   wire [1:0] _T_404 = _T_85 ? 2'h1 : _T_403; // @[Lookup.scala 34:39]
//   wire [1:0] _T_405 = _T_83 ? 2'h1 : _T_404; // @[Lookup.scala 34:39]
//   wire [1:0] _T_406 = _T_81 ? 2'h1 : _T_405; // @[Lookup.scala 34:39]
//   wire [1:0] _T_407 = _T_79 ? 2'h1 : _T_406; // @[Lookup.scala 34:39]
//   wire [1:0] _T_408 = _T_77 ? 2'h1 : _T_407; // @[Lookup.scala 34:39]
//   wire [1:0] _T_409 = _T_75 ? 2'h1 : _T_408; // @[Lookup.scala 34:39]
//   wire [1:0] _T_410 = _T_73 ? 2'h1 : _T_409; // @[Lookup.scala 34:39]
//   wire [1:0] _T_411 = _T_71 ? 2'h1 : _T_410; // @[Lookup.scala 34:39]
//   wire [1:0] _T_412 = _T_69 ? 2'h1 : _T_411; // @[Lookup.scala 34:39]
//   wire [1:0] _T_413 = _T_67 ? 2'h1 : _T_412; // @[Lookup.scala 34:39]
//   wire [1:0] _T_414 = _T_65 ? 2'h1 : _T_413; // @[Lookup.scala 34:39]
//   wire [1:0] _T_415 = _T_63 ? 2'h1 : _T_414; // @[Lookup.scala 34:39]
//   wire [1:0] _T_416 = _T_61 ? 2'h1 : _T_415; // @[Lookup.scala 34:39]
//   wire [1:0] _T_417 = _T_59 ? 2'h0 : _T_416; // @[Lookup.scala 34:39]
//   wire [1:0] _T_418 = _T_57 ? 2'h0 : _T_417; // @[Lookup.scala 34:39]
//   wire [1:0] _T_419 = _T_55 ? 2'h0 : _T_418; // @[Lookup.scala 34:39]
//   wire [1:0] _T_420 = _T_53 ? 2'h1 : _T_419; // @[Lookup.scala 34:39]
//   wire [1:0] _T_421 = _T_51 ? 2'h1 : _T_420; // @[Lookup.scala 34:39]
//   wire [1:0] _T_422 = _T_49 ? 2'h1 : _T_421; // @[Lookup.scala 34:39]
//   wire [1:0] _T_423 = _T_47 ? 2'h1 : _T_422; // @[Lookup.scala 34:39]
//   wire [1:0] _T_424 = _T_45 ? 2'h1 : _T_423; // @[Lookup.scala 34:39]
//   wire [1:0] _T_425 = _T_43 ? 2'h1 : _T_424; // @[Lookup.scala 34:39]
//   wire [1:0] _T_426 = _T_41 ? 2'h1 : _T_425; // @[Lookup.scala 34:39]
//   wire [1:0] _T_427 = _T_39 ? 2'h1 : _T_426; // @[Lookup.scala 34:39]
//   wire [1:0] _T_428 = _T_37 ? 2'h1 : _T_427; // @[Lookup.scala 34:39]
//   wire [1:0] _T_429 = _T_35 ? 2'h1 : _T_428; // @[Lookup.scala 34:39]
//   wire [1:0] _T_430 = _T_33 ? 2'h1 : _T_429; // @[Lookup.scala 34:39]
//   wire [1:0] _T_431 = _T_31 ? 2'h1 : _T_430; // @[Lookup.scala 34:39]
//   wire [1:0] _T_432 = _T_29 ? 2'h1 : _T_431; // @[Lookup.scala 34:39]
//   wire [1:0] _T_433 = _T_27 ? 2'h1 : _T_432; // @[Lookup.scala 34:39]
//   wire [1:0] _T_434 = _T_25 ? 2'h0 : _T_433; // @[Lookup.scala 34:39]
//   wire [1:0] _T_435 = _T_23 ? 2'h0 : _T_434; // @[Lookup.scala 34:39]
//   wire [1:0] _T_436 = _T_21 ? 2'h0 : _T_435; // @[Lookup.scala 34:39]
//   wire [1:0] _T_437 = _T_19 ? 2'h0 : _T_436; // @[Lookup.scala 34:39]
//   wire [1:0] _T_438 = _T_17 ? 2'h0 : _T_437; // @[Lookup.scala 34:39]
//   wire [1:0] _T_439 = _T_15 ? 2'h0 : _T_438; // @[Lookup.scala 34:39]
//   wire [1:0] _T_440 = _T_13 ? 2'h1 : _T_439; // @[Lookup.scala 34:39]
//   wire [1:0] _T_441 = _T_11 ? 2'h1 : _T_440; // @[Lookup.scala 34:39]
//   wire [1:0] _T_442 = _T_9 ? 2'h1 : _T_441; // @[Lookup.scala 34:39]
//   wire [1:0] _T_443 = _T_7 ? 2'h1 : _T_442; // @[Lookup.scala 34:39]
//   wire [1:0] _T_444 = _T_5 ? 2'h1 : _T_443; // @[Lookup.scala 34:39]
//   wire [1:0] _T_445 = _T_3 ? 2'h1 : _T_444; // @[Lookup.scala 34:39]
//   wire [1:0] dest_is_reg = _T_1 ? 2'h1 : _T_445; // @[Lookup.scala 34:39]
//   wire [1:0] _T_454 = _T_133 ? 2'h0 : _T_379; // @[Lookup.scala 34:39]
//   wire [1:0] _T_455 = _T_131 ? 2'h1 : _T_454; // @[Lookup.scala 34:39]
//   wire [1:0] _T_456 = _T_129 ? 2'h1 : _T_455; // @[Lookup.scala 34:39]
//   wire [1:0] _T_457 = _T_127 ? 2'h1 : _T_456; // @[Lookup.scala 34:39]
//   wire [1:0] _T_458 = _T_125 ? 2'h1 : _T_457; // @[Lookup.scala 34:39]
//   wire [1:0] _T_459 = _T_123 ? 2'h1 : _T_458; // @[Lookup.scala 34:39]
//   wire [1:0] _T_460 = _T_121 ? 2'h1 : _T_459; // @[Lookup.scala 34:39]
//   wire [1:0] _T_461 = _T_119 ? 2'h1 : _T_460; // @[Lookup.scala 34:39]
//   wire [1:0] _T_462 = _T_117 ? 2'h1 : _T_461; // @[Lookup.scala 34:39]
//   wire [1:0] _T_463 = _T_115 ? 2'h1 : _T_462; // @[Lookup.scala 34:39]
//   wire [1:0] _T_464 = _T_113 ? 2'h1 : _T_463; // @[Lookup.scala 34:39]
//   wire [1:0] _T_465 = _T_111 ? 2'h1 : _T_464; // @[Lookup.scala 34:39]
//   wire [1:0] _T_466 = _T_109 ? 2'h1 : _T_465; // @[Lookup.scala 34:39]
//   wire [1:0] _T_467 = _T_107 ? 2'h1 : _T_466; // @[Lookup.scala 34:39]
//   wire [1:0] _T_468 = _T_105 ? 2'h1 : _T_467; // @[Lookup.scala 34:39]
//   wire [1:0] _T_469 = _T_103 ? 2'h1 : _T_468; // @[Lookup.scala 34:39]
//   wire [1:0] _T_470 = _T_101 ? 2'h1 : _T_469; // @[Lookup.scala 34:39]
//   wire [1:0] _T_471 = _T_99 ? 2'h1 : _T_470; // @[Lookup.scala 34:39]
//   wire [1:0] _T_472 = _T_97 ? 2'h1 : _T_471; // @[Lookup.scala 34:39]
//   wire [1:0] _T_473 = _T_95 ? 2'h1 : _T_472; // @[Lookup.scala 34:39]
//   wire [1:0] _T_474 = _T_93 ? 2'h1 : _T_473; // @[Lookup.scala 34:39]
//   wire [1:0] _T_475 = _T_91 ? 2'h1 : _T_474; // @[Lookup.scala 34:39]
//   wire [1:0] _T_476 = _T_89 ? 2'h1 : _T_475; // @[Lookup.scala 34:39]
//   wire [1:0] _T_477 = _T_87 ? 2'h1 : _T_476; // @[Lookup.scala 34:39]
//   wire [1:0] _T_478 = _T_85 ? 2'h1 : _T_477; // @[Lookup.scala 34:39]
//   wire [1:0] _T_479 = _T_83 ? 2'h1 : _T_478; // @[Lookup.scala 34:39]
//   wire [1:0] _T_480 = _T_81 ? 2'h1 : _T_479; // @[Lookup.scala 34:39]
//   wire [1:0] _T_481 = _T_79 ? 2'h1 : _T_480; // @[Lookup.scala 34:39]
//   wire [1:0] _T_482 = _T_77 ? 2'h1 : _T_481; // @[Lookup.scala 34:39]
//   wire [1:0] _T_483 = _T_75 ? 2'h1 : _T_482; // @[Lookup.scala 34:39]
//   wire [1:0] _T_484 = _T_73 ? 2'h1 : _T_483; // @[Lookup.scala 34:39]
//   wire [1:0] _T_485 = _T_71 ? 2'h1 : _T_484; // @[Lookup.scala 34:39]
//   wire [1:0] _T_486 = _T_69 ? 2'h1 : _T_485; // @[Lookup.scala 34:39]
//   wire [1:0] _T_487 = _T_67 ? 2'h1 : _T_486; // @[Lookup.scala 34:39]
//   wire [1:0] _T_488 = _T_65 ? 2'h1 : _T_487; // @[Lookup.scala 34:39]
//   wire [1:0] _T_489 = _T_63 ? 2'h1 : _T_488; // @[Lookup.scala 34:39]
//   wire [1:0] _T_490 = _T_61 ? 2'h1 : _T_489; // @[Lookup.scala 34:39]
//   wire [1:0] _T_491 = _T_59 ? 2'h1 : _T_490; // @[Lookup.scala 34:39]
//   wire [1:0] _T_492 = _T_57 ? 2'h1 : _T_491; // @[Lookup.scala 34:39]
//   wire [1:0] _T_493 = _T_55 ? 2'h1 : _T_492; // @[Lookup.scala 34:39]
//   wire [1:0] _T_494 = _T_53 ? 2'h1 : _T_493; // @[Lookup.scala 34:39]
//   wire [1:0] _T_495 = _T_51 ? 2'h1 : _T_494; // @[Lookup.scala 34:39]
//   wire [1:0] _T_496 = _T_49 ? 2'h0 : _T_495; // @[Lookup.scala 34:39]
//   wire [1:0] _T_497 = _T_47 ? 2'h1 : _T_496; // @[Lookup.scala 34:39]
//   wire [1:0] _T_498 = _T_45 ? 2'h1 : _T_497; // @[Lookup.scala 34:39]
//   wire [1:0] _T_499 = _T_43 ? 2'h1 : _T_498; // @[Lookup.scala 34:39]
//   wire [1:0] _T_500 = _T_41 ? 2'h1 : _T_499; // @[Lookup.scala 34:39]
//   wire [1:0] _T_501 = _T_39 ? 2'h1 : _T_500; // @[Lookup.scala 34:39]
//   wire [1:0] _T_502 = _T_37 ? 2'h0 : _T_501; // @[Lookup.scala 34:39]
//   wire [1:0] _T_503 = _T_35 ? 2'h1 : _T_502; // @[Lookup.scala 34:39]
//   wire [1:0] _T_504 = _T_33 ? 2'h0 : _T_503; // @[Lookup.scala 34:39]
//   wire [1:0] _T_505 = _T_31 ? 2'h1 : _T_504; // @[Lookup.scala 34:39]
//   wire [1:0] _T_506 = _T_29 ? 2'h0 : _T_505; // @[Lookup.scala 34:39]
//   wire [1:0] _T_507 = _T_27 ? 2'h1 : _T_506; // @[Lookup.scala 34:39]
//   wire [1:0] _T_508 = _T_25 ? 2'h1 : _T_507; // @[Lookup.scala 34:39]
//   wire [1:0] _T_509 = _T_23 ? 2'h1 : _T_508; // @[Lookup.scala 34:39]
//   wire [1:0] _T_510 = _T_21 ? 2'h1 : _T_509; // @[Lookup.scala 34:39]
//   wire [1:0] _T_511 = _T_19 ? 2'h1 : _T_510; // @[Lookup.scala 34:39]
//   wire [1:0] _T_512 = _T_17 ? 2'h1 : _T_511; // @[Lookup.scala 34:39]
//   wire [1:0] _T_513 = _T_15 ? 2'h1 : _T_512; // @[Lookup.scala 34:39]
//   wire [1:0] _T_514 = _T_13 ? 2'h0 : _T_513; // @[Lookup.scala 34:39]
//   wire [1:0] _T_515 = _T_11 ? 2'h1 : _T_514; // @[Lookup.scala 34:39]
//   wire [1:0] _T_516 = _T_9 ? 2'h1 : _T_515; // @[Lookup.scala 34:39]
//   wire [1:0] _T_517 = _T_7 ? 2'h1 : _T_516; // @[Lookup.scala 34:39]
//   wire [1:0] _T_518 = _T_5 ? 2'h1 : _T_517; // @[Lookup.scala 34:39]
//   wire [1:0] _T_519 = _T_3 ? 2'h1 : _T_518; // @[Lookup.scala 34:39]
//   wire [1:0] rs1_is_reg = _T_1 ? 2'h1 : _T_519; // @[Lookup.scala 34:39]
//   wire [1:0] _T_529 = _T_131 ? 2'h1 : 2'h0; // @[Lookup.scala 34:39]
//   wire [1:0] _T_530 = _T_129 ? 2'h1 : _T_529; // @[Lookup.scala 34:39]
//   wire [1:0] _T_531 = _T_127 ? 2'h1 : _T_530; // @[Lookup.scala 34:39]
//   wire [1:0] _T_532 = _T_125 ? 2'h1 : _T_531; // @[Lookup.scala 34:39]
//   wire [1:0] _T_533 = _T_123 ? 2'h1 : _T_532; // @[Lookup.scala 34:39]
//   wire [1:0] _T_534 = _T_121 ? 2'h1 : _T_533; // @[Lookup.scala 34:39]
//   wire [1:0] _T_535 = _T_119 ? 2'h1 : _T_534; // @[Lookup.scala 34:39]
//   wire [1:0] _T_536 = _T_117 ? 2'h1 : _T_535; // @[Lookup.scala 34:39]
//   wire [1:0] _T_537 = _T_115 ? 2'h1 : _T_536; // @[Lookup.scala 34:39]
//   wire [1:0] _T_538 = _T_113 ? 2'h1 : _T_537; // @[Lookup.scala 34:39]
//   wire [1:0] _T_539 = _T_111 ? 2'h1 : _T_538; // @[Lookup.scala 34:39]
//   wire [1:0] _T_540 = _T_109 ? 2'h1 : _T_539; // @[Lookup.scala 34:39]
//   wire [1:0] _T_541 = _T_107 ? 2'h1 : _T_540; // @[Lookup.scala 34:39]
//   wire [1:0] _T_542 = _T_105 ? 2'h0 : _T_541; // @[Lookup.scala 34:39]
//   wire [1:0] _T_543 = _T_103 ? 2'h1 : _T_542; // @[Lookup.scala 34:39]
//   wire [1:0] _T_544 = _T_101 ? 2'h0 : _T_543; // @[Lookup.scala 34:39]
//   wire [1:0] _T_545 = _T_99 ? 2'h1 : _T_544; // @[Lookup.scala 34:39]
//   wire [1:0] _T_546 = _T_97 ? 2'h1 : _T_545; // @[Lookup.scala 34:39]
//   wire [1:0] _T_547 = _T_95 ? 2'h1 : _T_546; // @[Lookup.scala 34:39]
//   wire [1:0] _T_548 = _T_93 ? 2'h1 : _T_547; // @[Lookup.scala 34:39]
//   wire [1:0] _T_549 = _T_91 ? 2'h1 : _T_548; // @[Lookup.scala 34:39]
//   wire [1:0] _T_550 = _T_89 ? 2'h0 : _T_549; // @[Lookup.scala 34:39]
//   wire [1:0] _T_551 = _T_87 ? 2'h0 : _T_550; // @[Lookup.scala 34:39]
//   wire [1:0] _T_552 = _T_85 ? 2'h1 : _T_551; // @[Lookup.scala 34:39]
//   wire [1:0] _T_553 = _T_83 ? 2'h1 : _T_552; // @[Lookup.scala 34:39]
//   wire [1:0] _T_554 = _T_81 ? 2'h0 : _T_553; // @[Lookup.scala 34:39]
//   wire [1:0] _T_555 = _T_79 ? 2'h0 : _T_554; // @[Lookup.scala 34:39]
//   wire [1:0] _T_556 = _T_77 ? 2'h1 : _T_555; // @[Lookup.scala 34:39]
//   wire [1:0] _T_557 = _T_75 ? 2'h1 : _T_556; // @[Lookup.scala 34:39]
//   wire [1:0] _T_558 = _T_73 ? 2'h0 : _T_557; // @[Lookup.scala 34:39]
//   wire [1:0] _T_559 = _T_71 ? 2'h0 : _T_558; // @[Lookup.scala 34:39]
//   wire [1:0] _T_560 = _T_69 ? 2'h1 : _T_559; // @[Lookup.scala 34:39]
//   wire [1:0] _T_561 = _T_67 ? 2'h1 : _T_560; // @[Lookup.scala 34:39]
//   wire [1:0] _T_562 = _T_65 ? 2'h0 : _T_561; // @[Lookup.scala 34:39]
//   wire [1:0] _T_563 = _T_63 ? 2'h0 : _T_562; // @[Lookup.scala 34:39]
//   wire [1:0] _T_564 = _T_61 ? 2'h1 : _T_563; // @[Lookup.scala 34:39]
//   wire [1:0] _T_565 = _T_59 ? 2'h1 : _T_564; // @[Lookup.scala 34:39]
//   wire [1:0] _T_566 = _T_57 ? 2'h1 : _T_565; // @[Lookup.scala 34:39]
//   wire [1:0] _T_567 = _T_55 ? 2'h1 : _T_566; // @[Lookup.scala 34:39]
//   wire [1:0] _T_568 = _T_53 ? 2'h0 : _T_567; // @[Lookup.scala 34:39]
//   wire [1:0] _T_569 = _T_51 ? 2'h0 : _T_568; // @[Lookup.scala 34:39]
//   wire [1:0] _T_570 = _T_49 ? 2'h0 : _T_569; // @[Lookup.scala 34:39]
//   wire [1:0] _T_571 = _T_47 ? 2'h0 : _T_570; // @[Lookup.scala 34:39]
//   wire [1:0] _T_572 = _T_45 ? 2'h0 : _T_571; // @[Lookup.scala 34:39]
//   wire [1:0] _T_573 = _T_43 ? 2'h0 : _T_572; // @[Lookup.scala 34:39]
//   wire [1:0] _T_574 = _T_41 ? 2'h0 : _T_573; // @[Lookup.scala 34:39]
//   wire [1:0] _T_575 = _T_39 ? 2'h0 : _T_574; // @[Lookup.scala 34:39]
//   wire [1:0] _T_576 = _T_37 ? 2'h0 : _T_575; // @[Lookup.scala 34:39]
//   wire [1:0] _T_577 = _T_35 ? 2'h0 : _T_576; // @[Lookup.scala 34:39]
//   wire [1:0] _T_578 = _T_33 ? 2'h0 : _T_577; // @[Lookup.scala 34:39]
//   wire [1:0] _T_579 = _T_31 ? 2'h0 : _T_578; // @[Lookup.scala 34:39]
//   wire [1:0] _T_580 = _T_29 ? 2'h0 : _T_579; // @[Lookup.scala 34:39]
//   wire [1:0] _T_581 = _T_27 ? 2'h0 : _T_580; // @[Lookup.scala 34:39]
//   wire [1:0] _T_582 = _T_25 ? 2'h1 : _T_581; // @[Lookup.scala 34:39]
//   wire [1:0] _T_583 = _T_23 ? 2'h1 : _T_582; // @[Lookup.scala 34:39]
//   wire [1:0] _T_584 = _T_21 ? 2'h1 : _T_583; // @[Lookup.scala 34:39]
//   wire [1:0] _T_585 = _T_19 ? 2'h1 : _T_584; // @[Lookup.scala 34:39]
//   wire [1:0] _T_586 = _T_17 ? 2'h1 : _T_585; // @[Lookup.scala 34:39]
//   wire [1:0] _T_587 = _T_15 ? 2'h1 : _T_586; // @[Lookup.scala 34:39]
//   wire [1:0] _T_588 = _T_13 ? 2'h0 : _T_587; // @[Lookup.scala 34:39]
//   wire [1:0] _T_589 = _T_11 ? 2'h0 : _T_588; // @[Lookup.scala 34:39]
//   wire [1:0] _T_590 = _T_9 ? 2'h1 : _T_589; // @[Lookup.scala 34:39]
//   wire [1:0] _T_591 = _T_7 ? 2'h1 : _T_590; // @[Lookup.scala 34:39]
//   wire [1:0] _T_592 = _T_5 ? 2'h0 : _T_591; // @[Lookup.scala 34:39]
//   wire [1:0] _T_593 = _T_3 ? 2'h0 : _T_592; // @[Lookup.scala 34:39]
//   wire [1:0] rs2_is_reg = _T_1 ? 2'h1 : _T_593; // @[Lookup.scala 34:39]
//   wire [19:0] _imm_data_T_2 = io_get_inst_bits_inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 77:12]
//   wire [31:0] _imm_data_T_4 = {_imm_data_T_2,csr_addr}; // @[Cat.scala 33:92]
//   wire [31:0] _imm_data_T_6 = {io_get_inst_bits_inst[31:12],12'h0}; // @[Cat.scala 33:92]
//   wire [31:0] _imm_data_T_13 = {_imm_data_T_2,io_get_inst_bits_inst[31:25],dest_addr}; // @[Cat.scala 33:92]
//   wire [11:0] _imm_data_T_16 = io_get_inst_bits_inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 77:12]
//   wire [31:0] _imm_data_T_23 = {_imm_data_T_16,io_get_inst_bits_inst[19:12],io_get_inst_bits_inst[20],
//     io_get_inst_bits_inst[30:21],1'h0}; // @[Cat.scala 33:92]
//   wire [31:0] _imm_data_T_33 = {_imm_data_T_2,io_get_inst_bits_inst[7],io_get_inst_bits_inst[30:25],
//     io_get_inst_bits_inst[11:8],1'h0}; // @[Cat.scala 33:92]
//   wire [31:0] _imm_data_T_35 = {27'h0,rs1_addr}; // @[Cat.scala 33:92]
//   wire [31:0] _imm_data_T_37 = {26'h0,io_get_inst_bits_inst[25:20]}; // @[Cat.scala 33:92]
//   wire [31:0] _imm_data_T_39 = 4'hc == instType ? _imm_data_T_4 : 32'h0; // @[Mux.scala 81:58]
//   wire [31:0] _imm_data_T_41 = 4'h1 == instType ? _imm_data_T_6 : _imm_data_T_39; // @[Mux.scala 81:58]
//   wire [31:0] _imm_data_T_43 = 4'h3 == instType ? _imm_data_T_13 : _imm_data_T_41; // @[Mux.scala 81:58]
//   wire [31:0] _imm_data_T_45 = 4'h2 == instType ? _imm_data_T_23 : _imm_data_T_43; // @[Mux.scala 81:58]
//   wire [31:0] _imm_data_T_47 = 4'h7 == instType ? _imm_data_T_33 : _imm_data_T_45; // @[Mux.scala 81:58]
//   wire  temp_rs1_is_reg = rs1_is_reg == 2'h1; // @[decode.scala 73:43]
//   wire  temp_rs2_is_reg = rs2_is_reg == 2'h1; // @[decode.scala 74:43]
//   wire [1:0] _GEN_12 = io_op_datas_ready ? dest_is_reg : {{1'd0}, reg_dest_is_reg}; // @[decode.scala 79:20 94:33 42:38]
//   wire [1:0] _GEN_16 = reset ? 2'h0 : _GEN_12; // @[decode.scala 42:{38,38}]
//   assign io_get_inst_ready = io_op_datas_ready; // @[decode.scala 21:31]
//   assign io_normal_rd_rs1_addr = io_get_inst_bits_inst[19:15]; // @[decode.scala 55:35]
//   assign io_normal_rd_rs2_addr = io_get_inst_bits_inst[24:20]; // @[decode.scala 54:35]
//   assign io_csr_rd_csr_addr = io_get_inst_bits_inst[31:20]; // @[decode.scala 56:35]
//   assign io_op_datas_valid = reg_valid; // @[decode.scala 120:57]
//   assign io_op_datas_bits_opType = reg_opType; // @[decode.scala 105:49]
//   assign io_op_datas_bits_exuType = reg_exuType; // @[decode.scala 106:49]
//   assign io_op_datas_bits_rs1_addr = reg_rs1_addr; // @[decode.scala 107:49]
//   assign io_op_datas_bits_rs1_data = reg_rs1_data; // @[decode.scala 108:49]
//   assign io_op_datas_bits_rs2_addr = reg_rs2_addr; // @[decode.scala 109:49]
//   assign io_op_datas_bits_rs2_data = reg_rs2_data; // @[decode.scala 110:49]
//   assign io_op_datas_bits_imm = reg_imm; // @[decode.scala 111:49]
//   assign io_op_datas_bits_pc = reg_pc; // @[decode.scala 112:57]
//   assign io_op_datas_bits_inst = reg_inst; // @[decode.scala 113:49]
//   assign io_op_datas_bits_dest_addr = reg_dest_addr; // @[decode.scala 114:49]
//   assign io_op_datas_bits_dest_is_reg = reg_dest_is_reg; // @[decode.scala 115:41]
//   assign io_op_datas_bits_is_pre = reg_is_pre; // @[decode.scala 119:49]
//   assign io_op_datas_bits_csr_addr = reg_csr_addr; // @[decode.scala 117:49]
//   assign io_op_datas_bits_csr_data = reg_csr_data; // @[decode.scala 118:49]

// always @(posedge clock)begin 
// 	if(reset)begin 
// 		reg_valid <= 1'h0;
// 	end else if (io_flush) begin 
// 		reg_valid <= 1'h0;
// 	end else if (io_op_datas_ready) begin
// 		reg_valid <= io_get_inst_valid;
// 	end 
// end

// always @(posedge clock)begin 
// 	if(reset)begin 
// 		reg_opType <= 3'h0;
// 		reg_exuType <= 7'h0;
// 		reg_rs1_addr <= 5'h0;
// 		reg_rs1_data <= 64'h0;
// 		reg_rs2_addr <= 5'h0;
// 		reg_rs2_data <= 64'h0;
// 		reg_imm <= 32'h0;
// 		reg_pc <= 64'h0;
// 		reg_inst <= 32'h0;
// 		reg_dest_addr <= 5'h0;
// 		reg_csr_addr <= 12'h0;
// 		reg_csr_data <= 64'h0;
// 		reg_is_pre <= 1'h0;
// 	end else if(io_op_datas_ready)begin 
//       if (_T_1) begin // @[Lookup.scala 34:39]
//         reg_opType <= 3'h2;
// 		reg_exuType <= 7'h2;
//       end else if (_T_3) begin // @[Lookup.scala 34:39]
//         reg_opType <= 3'h2;
// 		reg_exuType <= 7'h0;
//       end else begin
//         reg_opType <= _T_222;
// 		reg_exuType <= _T_296;
//       end
//       if (temp_rs1_is_reg) begin // @[decode.scala 75:34]
//         reg_rs1_addr <= rs1_addr;
// 		reg_rs1_data <= io_normal_rd_rs1_data;
//       end else begin
//         reg_rs1_addr <= 5'h0;
// 		reg_rs1_data <= 64'h0;
//       end
//       if (temp_rs2_is_reg) begin // @[decode.scala 77:34]
//         reg_rs2_addr <= rs2_addr;
// 		reg_rs2_data <= io_normal_rd_rs2_data;
//       end else begin
//         reg_rs2_addr <= 5'h0;
// 		reg_rs2_data <= 64'h0;
//       end

//       if (4'h4 == instType) begin // @[Mux.scala 81:58]
//         reg_imm <= _imm_data_T_37;
//       end else if (4'h5 == instType) begin // @[Mux.scala 81:58]
//         reg_imm <= _imm_data_T_35;
//       end else begin
//         reg_imm <= _imm_data_T_47;
//       end
// 	  reg_pc <= io_get_inst_bits_pc;
// 	  reg_inst <= io_get_inst_bits_inst;
// 	  reg_dest_addr <= dest_addr;
// 	  reg_csr_addr <= csr_addr;
// 	  reg_csr_data <= io_csr_rd_csr_data;
// 	  reg_is_pre <= io_get_inst_bits_is_pre;
// 	end
// 	reg_dest_is_reg <= _GEN_16[0];
// end 
endmodule